-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition
-- Created on Mon Sep 24 20:43:10 2018

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM1 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        input1 : IN STD_LOGIC := '0';
        output1 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
    );
END SM1;

ARCHITECTURE BEHAVIOR OF SM1 IS
    TYPE type_fstate IS (state1,state4,state7,state10,state5,state3,state2,state6,state8,state9,state11,state14,state13,state15,state12,state16,state17,state18);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,input1)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            output1 <= "00000000000000";
        ELSE
            output1 <= "00000000000000";
            CASE fstate IS
                WHEN state1 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    output1 <= "00100001000000";
                WHEN state4 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    output1 <= "00100100100000";
                WHEN state7 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;

                    output1 <= "00101000010000";
                WHEN state10 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state11;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state10;
                    END IF;

                    output1 <= "00101100001000";
                WHEN state5 =>
                    IF (NOT((input1 = '1'))) THEN
                        reg_fstate <= state4;
                    ELSIF ((input1 = '1')) THEN
                        reg_fstate <= state6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    output1 <= "10000110000000";
                WHEN state3 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    output1 <= "00000011000000";
                WHEN state2 =>
                    IF (NOT((input1 = '1'))) THEN
                        reg_fstate <= state1;
                    ELSIF ((input1 = '1')) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    output1 <= "10100010000000";
                WHEN state6 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;

                    output1 <= "00000110100000";
                WHEN state8 =>
                    IF (NOT((input1 = '1'))) THEN
                        reg_fstate <= state7;
                    ELSIF ((input1 = '1')) THEN
                        reg_fstate <= state9;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state8;
                    END IF;

                    output1 <= "10101010000000";
                WHEN state9 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state9;
                    END IF;

                    output1 <= "00001010010000";
                WHEN state11 =>
                    IF (NOT((input1 = '1'))) THEN
                        reg_fstate <= state10;
                    ELSIF ((input1 = '1')) THEN
                        reg_fstate <= state12;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state11;
                    END IF;

                    output1 <= "10001110000000";
                WHEN state14 =>
                    IF (NOT((input1 = '1'))) THEN
                        reg_fstate <= state13;
                    ELSIF ((input1 = '1')) THEN
                        reg_fstate <= state15;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state14;
                    END IF;

                    output1 <= "01110010000000";
                WHEN state13 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state14;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state13;
                    END IF;

                    output1 <= "00110000000100";
                WHEN state15 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state16;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state15;
                    END IF;

                    output1 <= "00010010000100";
                WHEN state12 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state13;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state12;
                    END IF;

                    output1 <= "00001110001000";
                WHEN state16 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state17;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state16;
                    END IF;

                    output1 <= "00110100000010";
                WHEN state17 =>
                    IF (NOT((input1 = '1'))) THEN
                        reg_fstate <= state16;
                    ELSIF ((input1 = '1')) THEN
                        reg_fstate <= state18;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state17;
                    END IF;

                    output1 <= "01010110000000";
                WHEN state18 =>
                    IF ((input1 = '1')) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state18;
                    END IF;

                    output1 <= "00010110000010";
                WHEN OTHERS => 
                    output1 <= "XXXXXXXXXXXXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
